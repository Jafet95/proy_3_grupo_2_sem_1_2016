`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: Jafet Chaves Barrantes
// 
// Create Date:    21:04:45 05/26/2016 
// Design Name: 
// Module Name:    prueba_lectura_rtc 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module prueba_lectura_rtc(
    );
//Aqu� va la instanciaci�n del microcontrolador, el banco de registros y el control con la
//respectiva interfaz con el PicoBlaze
//No hace falta el Demux como el proyecto pasado

endmodule
